class adder_transaction;
    logic [3:0] op_a;
    logic [3:0] op_b;
    logic carry_in;
    logic [3:0] sum;
    logic carry_out;

    // function void display(string name);
    //     $display("-------------------------");
    //     $display("- %s ",name);
    //     $display("-------------------------");
    //     $display("- a = %0d, b = %0d",a,b);
    //     $display("- c = %0d",c);
    //     $display("-------------------------");
    // endfunction 
endclass