interface adder_intf();
    bit [3:0] op_a;
    bit [3:0] op_b;
    bit carry_in;
    bit [3:0] sum;
    bit carry_out;
endinterface
