interface adder_intf();
    logic [3:0] op_a;
    logic [3:0] op_b;
    logic carry_in;
    logic [3:0] sum;
    logic carry_out;
endinterface
